module hadder
{
input a,b
output sum,carry
};
sum=a^b;
carry=a&b;
endmodule 
